module Instr_Mem(input logic[7:0] A, output logic[31:0] RD);
	always_comb begin
		case(A)
			8'b00000000: RD = 32'b_001000_00000_00001_00000_00011_001010;
			8'b00000001: RD = 32'b_000000_00001_00001_00001_00000_100000;
			8'b00000010: RD = 32'b_000000_00001_00001_00001_00000_100000;
			8'b00000011: RD = 32'b_000000_00001_00001_00001_00000_100000;
			8'b00000100: RD = 32'b_000000_00001_00001_00001_00000_100000;
			8'b00000101: RD = 32'b_000000_00001_00010_00101_00000_100111;
			8'b00000110: RD = 32'b_000000_00101_00100_00110_00000_101010;
			default: RD = 32'b_000000_00000_00000_00000_00000_000000;
		endcase
	end
endmodule 